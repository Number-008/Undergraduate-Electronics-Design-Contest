library verilog;
use verilog.vl_types.all;
entity DDS_vlg_tst is
end DDS_vlg_tst;
